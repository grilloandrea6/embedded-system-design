module rgb565Grayscalelse #(parameter [7:0] customInstructionId = 8'd0)
                (input wire start,
                input wire [31:0] valueA,
                input wire [7:0] isId,
                output wire done,
                output wire [31:0] result);



endmodule